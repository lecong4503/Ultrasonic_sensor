`timescale 1ns / 1ps

module echo (
    input clk,
    input rst_n,
    input us_cnt,
    input ms_cnt,
    
)